
module nios (
	clk_clk,
	reset_reset_n,
	gpio_out_external_connection_export,
	switch_external_connection_export);	

	input		clk_clk;
	input		reset_reset_n;
	output		gpio_out_external_connection_export;
	input		switch_external_connection_export;
endmodule
